module top(//8-3优先编码器
    input [7:0] x,
    input en,
    output reg p,
    output reg [2:0] y,
    output reg [7:0] HEX
);
    wire [3:0] yh;
    always @(*)begin
        if(en)begin
            p = 1'b0;
            y = 3'b000;
            for(integer i=0;i<=7;i=i+1)begin
                if(x[i]==1'b1) begin
                    y = i[2:0];
                    p = 1'b1;
                end
            end
        end
        else begin
            y=3'b000;
            p=1'b0;
        end
        if(y==3'b000)begin
            p = 1'b0;
        end
    end
    assign yh = en?{1'b0,y}:4'b1111;
    bcd7seg bcd7seg_moudle(
        .b(yh),
        .h(HEX[7:0])
    );
endmodule

module bcd7seg(
    input [3:0] b,
    output reg [7:0] h
);
always @(*)begin
    case(b)
        4'b0000 : h = 8'b00000011;
        4'b0001 : h = 8'b10011111;
        4'b0010 : h = 8'b00100101;
        4'b0011 : h = 8'b00001101;
        4'b0100 : h = 8'b10011001;
        4'b0101 : h = 8'b01001001;
        4'b0110 : h = 8'b01000001;
        4'b0111 : h = 8'b00011111;
        4'b1000 : h = 8'b00000001;
        4'b1001 : h = 8'b00001001;
        default: h = 8'b11111111;
    endcase
end
endmodule